* SPICE NETLIST
***************************************

.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_2t PLUS MINUS
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT fmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT fmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lincap PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lincap_rf_25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lowcpad_d15 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d23 APAD AVSS
.ENDS
***************************************
.SUBCKT mimcap_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ndio_hia_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwod D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_cas_nw D GB S B GT
.ENDS
***************************************
.SUBCKT nmos_rf_cross_nw DP DM S B
.ENDS
***************************************
.SUBCKT nmos_rf_diff_nw DP GP S B DM GM
.ENDS
***************************************
.SUBCKT nmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_na18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_rdk D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_lpg PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_hia_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwod D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_rdk D G S B
.ENDS
***************************************
.SUBCKT pmoscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT probe1 TOP BULK
.ENDS
***************************************
.SUBCKT probe2 TOP BULK
.ENDS
***************************************
.SUBCKT probe3 TOP BULK
.ENDS
***************************************
.SUBCKT probe4 TOP BULK
.ENDS
***************************************
.SUBCKT probe5 TOP BULK
.ENDS
***************************************
.SUBCKT probe6 TOP BULK
.ENDS
***************************************
.SUBCKT probe7 TOP BULK
.ENDS
***************************************
.SUBCKT rfesd_rf1 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf2 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf3 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf4 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf5 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf6 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf7 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf8 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sline_gscpw_mu PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sline_ms_mu PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z_rdk PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT TAPCELLBWP7T
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT DFCNQD1BWP7T CP D CDN VDD VSS Q
** N=19 EP=6 IP=0 FDC=28
M0 VSS CP 7 VSS nch L=6e-08 W=1.5e-07 $X=230 $Y=200 $D=4
M1 9 7 VSS VSS nch L=6e-08 W=1.5e-07 $X=520 $Y=345 $D=4
M2 16 7 VSS VSS nch L=6e-08 W=1.6e-07 $X=980 $Y=240 $D=4
M3 8 D 16 VSS nch L=6e-08 W=1.6e-07 $X=1170 $Y=240 $D=4
M4 17 9 8 VSS nch L=6e-08 W=1.5e-07 $X=1505 $Y=350 $D=4
M5 18 10 17 VSS nch L=6e-08 W=1.5e-07 $X=1755 $Y=220 $D=4
M6 VSS CDN 18 VSS nch L=6e-08 W=1.5e-07 $X=1955 $Y=220 $D=4
M7 10 8 VSS VSS nch L=6e-08 W=1.5e-07 $X=2315 $Y=200 $D=4
M8 12 9 10 VSS nch L=6e-08 W=1.5e-07 $X=2660 $Y=350 $D=4
M9 11 7 12 VSS nch L=6e-08 W=1.5e-07 $X=2950 $Y=400 $D=4
M10 VSS 13 11 VSS nch L=6e-08 W=1.5e-07 $X=3500 $Y=220 $D=4
M11 19 CDN VSS VSS nch L=6e-08 W=3e-07 $X=3810 $Y=235 $D=4
M12 13 12 19 VSS nch L=6e-08 W=3e-07 $X=4010 $Y=235 $D=4
M13 Q 13 VSS VSS nch L=6e-08 W=3e-07 $X=4500 $Y=200 $D=4
M14 VDD CP 7 VDD pch L=6e-08 W=1.9e-07 $X=230 $Y=820 $D=103
M15 9 7 VDD VDD pch L=6e-08 W=1.7e-07 $X=470 $Y=820 $D=103
M16 14 9 VDD VDD pch L=6e-08 W=1.6e-07 $X=960 $Y=820 $D=103
M17 8 D 14 VDD pch L=6e-08 W=1.6e-07 $X=1150 $Y=820 $D=103
M18 15 7 8 VDD pch L=6e-08 W=1.5e-07 $X=1470 $Y=900 $D=103
M19 VDD 10 15 VDD pch L=6e-08 W=1.5e-07 $X=1710 $Y=900 $D=103
M20 VDD CDN 15 VDD pch L=6e-08 W=1.5e-07 $X=2200 $Y=1030 $D=103
M21 10 8 VDD VDD pch L=6e-08 W=1.5e-07 $X=2520 $Y=870 $D=103
M22 12 7 10 VDD pch L=6e-08 W=1.5e-07 $X=2875 $Y=870 $D=103
M23 11 9 12 VDD pch L=6e-08 W=1.5e-07 $X=3200 $Y=870 $D=103
M24 VDD 13 11 VDD pch L=6e-08 W=1.5e-07 $X=3460 $Y=870 $D=103
M25 13 CDN VDD VDD pch L=6e-08 W=1.9e-07 $X=3830 $Y=985 $D=103
M26 VDD 12 13 VDD pch L=6e-08 W=3.2e-07 $X=4090 $Y=855 $D=103
M27 Q 13 VDD VDD pch L=6e-08 W=3.45e-07 $X=4500 $Y=855 $D=103
.ENDS
***************************************
.SUBCKT lfsr4
** N=34 EP=0 IP=22 FDC=134
M0 22 1 2 22 nch L=6e-08 W=1.5e-07 $X=4060 $Y=1565 $D=4
M1 3 2 22 22 nch L=6e-08 W=3e-07 $X=4340 $Y=1565 $D=4
M2 22 3 4 22 nch L=6e-08 W=1.2e-07 $X=4875 $Y=1580 $D=4
M3 5 4 22 22 nch L=6e-08 W=1.2e-07 $X=5135 $Y=1580 $D=4
M4 6 5 22 22 nch L=6e-08 W=1.5e-07 $X=5760 $Y=1565 $D=4
M5 22 7 8 22 nch L=6e-08 W=3e-07 $X=6250 $Y=1565 $D=4
M6 30 9 22 22 nch L=6e-08 W=1.5e-07 $X=6520 $Y=1765 $D=4
M7 11 7 30 22 nch L=6e-08 W=1.5e-07 $X=6780 $Y=1595 $D=4
M8 9 8 11 22 nch L=6e-08 W=1.8e-07 $X=7040 $Y=1565 $D=4
M9 22 10 9 22 nch L=6e-08 W=1.8e-07 $X=7390 $Y=1685 $D=4
M10 12 11 22 22 nch L=6e-08 W=1.95e-07 $X=7750 $Y=1670 $D=4
M11 22 13 16 22 nch L=6e-08 W=1.5e-07 $X=8260 $Y=1715 $D=4
M12 15 16 22 22 nch L=6e-08 W=1.5e-07 $X=8500 $Y=1715 $D=4
M13 31 16 22 22 nch L=6e-08 W=2.8e-07 $X=8960 $Y=1585 $D=4
M14 17 14 31 22 nch L=6e-08 W=2.8e-07 $X=9160 $Y=1585 $D=4
M15 32 15 17 22 nch L=6e-08 W=1.5e-07 $X=9430 $Y=1715 $D=4
M16 22 18 32 22 nch L=6e-08 W=1.5e-07 $X=9705 $Y=1745 $D=4
M17 33 17 22 22 nch L=6e-08 W=1.5e-07 $X=10085 $Y=1745 $D=4
M18 18 6 33 22 nch L=6e-08 W=1.5e-07 $X=10285 $Y=1745 $D=4
M19 20 15 18 22 nch L=6e-08 W=1.5e-07 $X=10545 $Y=1745 $D=4
M20 19 16 20 22 nch L=6e-08 W=1.5e-07 $X=10805 $Y=1745 $D=4
M21 34 6 19 22 nch L=6e-08 W=1.5e-07 $X=11345 $Y=1745 $D=4
M22 22 21 34 22 nch L=6e-08 W=1.5e-07 $X=11560 $Y=1745 $D=4
M23 21 20 22 22 nch L=6e-08 W=3.1e-07 $X=11900 $Y=1585 $D=4
M24 24 21 22 22 nch L=6e-08 W=2.8e-07 $X=12485 $Y=1585 $D=4
M25 23 1 2 23 pch L=6e-08 W=1.9e-07 $X=4060 $Y=2375 $D=103
M26 3 2 23 23 pch L=6e-08 W=3.8e-07 $X=4340 $Y=2185 $D=103
M27 23 3 4 23 pch L=6e-08 W=2.25e-07 $X=4860 $Y=2340 $D=103
M28 5 4 23 23 pch L=6e-08 W=2.25e-07 $X=5120 $Y=2340 $D=103
M29 6 5 23 23 pch L=6e-08 W=1.9e-07 $X=5760 $Y=2375 $D=103
M30 23 7 8 23 pch L=6e-08 W=1.5e-07 $X=6250 $Y=2415 $D=103
M31 27 9 23 23 pch L=6e-08 W=1.5e-07 $X=6585 $Y=2235 $D=103
M32 11 8 27 23 pch L=6e-08 W=1.5e-07 $X=6800 $Y=2235 $D=103
M33 9 7 11 23 pch L=6e-08 W=1.5e-07 $X=7140 $Y=2415 $D=103
M34 23 10 9 23 pch L=6e-08 W=1.9e-07 $X=7400 $Y=2375 $D=103
M35 12 11 23 23 pch L=6e-08 W=1.5e-07 $X=7750 $Y=2415 $D=103
M36 23 13 16 23 pch L=6e-08 W=1.9e-07 $X=8260 $Y=2185 $D=103
M37 15 16 23 23 pch L=6e-08 W=1.9e-07 $X=8500 $Y=2185 $D=103
M38 28 15 23 23 pch L=6e-08 W=1.9e-07 $X=9015 $Y=2335 $D=103
M39 17 14 28 23 pch L=6e-08 W=1.9e-07 $X=9205 $Y=2335 $D=103
M40 29 16 17 23 pch L=6e-08 W=1.5e-07 $X=9490 $Y=2265 $D=103
M41 23 18 29 23 pch L=6e-08 W=1.5e-07 $X=9765 $Y=2215 $D=103
M42 18 17 23 23 pch L=6e-08 W=1.5e-07 $X=10045 $Y=2215 $D=103
M43 23 6 18 23 pch L=6e-08 W=1.5e-07 $X=10305 $Y=2215 $D=103
M44 20 16 18 23 pch L=6e-08 W=1.5e-07 $X=10780 $Y=2215 $D=103
M45 19 15 20 23 pch L=6e-08 W=1.5e-07 $X=11040 $Y=2215 $D=103
M46 23 6 19 23 pch L=6e-08 W=1.95e-07 $X=11300 $Y=2215 $D=103
M47 19 21 23 23 pch L=6e-08 W=1.6e-07 $X=11540 $Y=2215 $D=103
M48 21 20 23 23 pch L=6e-08 W=3.25e-07 $X=12015 $Y=2220 $D=103
M49 24 21 23 23 pch L=6e-08 W=3.8e-07 $X=12525 $Y=2185 $D=103
X52 13 24 6 23 22 25 DFCNQD1BWP7T $T=12835 1365 0 0 $X=12600 $Y=1260
X53 13 25 6 23 22 7 DFCNQD1BWP7T $T=17635 1365 0 0 $X=17400 $Y=1260
X54 26 7 6 23 22 10 DFCNQD1BWP7T $T=22435 1365 0 0 $X=22200 $Y=1260
.ENDS
***************************************
